// AND Gate
module and2(x,y,s);
input x,y;
output s;

//2. RTL M
assign s=x&y;

endmodule
